module gamma(input [7:0] in, output [11:0] out);
assign out =  	(in == 8'h00) ? 12'h000 : 
	(in == 8'h01) ? 12'h000 : 
	(in == 8'h02) ? 12'h000 : 
	(in == 8'h03) ? 12'h001 : 
	(in == 8'h04) ? 12'h001 : 
	(in == 8'h05) ? 12'h002 : 
	(in == 8'h06) ? 12'h002 : 
	(in == 8'h07) ? 12'h003 : 
	(in == 8'h08) ? 12'h004 : 
	(in == 8'h09) ? 12'h005 : 
	(in == 8'h0a) ? 12'h006 : 
	(in == 8'h0b) ? 12'h008 : 
	(in == 8'h0c) ? 12'h009 : 
	(in == 8'h0d) ? 12'h00b : 
	(in == 8'h0e) ? 12'h00c : 
	(in == 8'h0f) ? 12'h00e : 
	(in == 8'h10) ? 12'h010 : 
	(in == 8'h11) ? 12'h012 : 
	(in == 8'h12) ? 12'h014 : 
	(in == 8'h13) ? 12'h017 : 
	(in == 8'h14) ? 12'h019 : 
	(in == 8'h15) ? 12'h01c : 
	(in == 8'h16) ? 12'h01e : 
	(in == 8'h17) ? 12'h021 : 
	(in == 8'h18) ? 12'h024 : 
	(in == 8'h19) ? 12'h027 : 
	(in == 8'h1a) ? 12'h02b : 
	(in == 8'h1b) ? 12'h02e : 
	(in == 8'h1c) ? 12'h031 : 
	(in == 8'h1d) ? 12'h035 : 
	(in == 8'h1e) ? 12'h039 : 
	(in == 8'h1f) ? 12'h03d : 
	(in == 8'h20) ? 12'h040 : 
	(in == 8'h21) ? 12'h045 : 
	(in == 8'h22) ? 12'h049 : 
	(in == 8'h23) ? 12'h04d : 
	(in == 8'h24) ? 12'h052 : 
	(in == 8'h25) ? 12'h056 : 
	(in == 8'h26) ? 12'h05b : 
	(in == 8'h27) ? 12'h060 : 
	(in == 8'h28) ? 12'h065 : 
	(in == 8'h29) ? 12'h06a : 
	(in == 8'h2a) ? 12'h06f : 
	(in == 8'h2b) ? 12'h074 : 
	(in == 8'h2c) ? 12'h07a : 
	(in == 8'h2d) ? 12'h080 : 
	(in == 8'h2e) ? 12'h085 : 
	(in == 8'h2f) ? 12'h08b : 
	(in == 8'h30) ? 12'h091 : 
	(in == 8'h31) ? 12'h097 : 
	(in == 8'h32) ? 12'h09d : 
	(in == 8'h33) ? 12'h0a4 : 
	(in == 8'h34) ? 12'h0aa : 
	(in == 8'h35) ? 12'h0b1 : 
	(in == 8'h36) ? 12'h0b8 : 
	(in == 8'h37) ? 12'h0bf : 
	(in == 8'h38) ? 12'h0c5 : 
	(in == 8'h39) ? 12'h0cd : 
	(in == 8'h3a) ? 12'h0d4 : 
	(in == 8'h3b) ? 12'h0db : 
	(in == 8'h3c) ? 12'h0e3 : 
	(in == 8'h3d) ? 12'h0ea : 
	(in == 8'h3e) ? 12'h0f2 : 
	(in == 8'h3f) ? 12'h0fa : 
	(in == 8'h40) ? 12'h102 : 
	(in == 8'h41) ? 12'h10a : 
	(in == 8'h42) ? 12'h112 : 
	(in == 8'h43) ? 12'h11b : 
	(in == 8'h44) ? 12'h123 : 
	(in == 8'h45) ? 12'h12c : 
	(in == 8'h46) ? 12'h135 : 
	(in == 8'h47) ? 12'h13d : 
	(in == 8'h48) ? 12'h146 : 
	(in == 8'h49) ? 12'h150 : 
	(in == 8'h4a) ? 12'h159 : 
	(in == 8'h4b) ? 12'h162 : 
	(in == 8'h4c) ? 12'h16c : 
	(in == 8'h4d) ? 12'h175 : 
	(in == 8'h4e) ? 12'h17f : 
	(in == 8'h4f) ? 12'h189 : 
	(in == 8'h50) ? 12'h193 : 
	(in == 8'h51) ? 12'h19d : 
	(in == 8'h52) ? 12'h1a7 : 
	(in == 8'h53) ? 12'h1b2 : 
	(in == 8'h54) ? 12'h1bc : 
	(in == 8'h55) ? 12'h1c7 : 
	(in == 8'h56) ? 12'h1d2 : 
	(in == 8'h57) ? 12'h1dd : 
	(in == 8'h58) ? 12'h1e8 : 
	(in == 8'h59) ? 12'h1f3 : 
	(in == 8'h5a) ? 12'h1fe : 
	(in == 8'h5b) ? 12'h20a : 
	(in == 8'h5c) ? 12'h215 : 
	(in == 8'h5d) ? 12'h221 : 
	(in == 8'h5e) ? 12'h22c : 
	(in == 8'h5f) ? 12'h238 : 
	(in == 8'h60) ? 12'h244 : 
	(in == 8'h61) ? 12'h251 : 
	(in == 8'h62) ? 12'h25d : 
	(in == 8'h63) ? 12'h269 : 
	(in == 8'h64) ? 12'h276 : 
	(in == 8'h65) ? 12'h282 : 
	(in == 8'h66) ? 12'h28f : 
	(in == 8'h67) ? 12'h29c : 
	(in == 8'h68) ? 12'h2a9 : 
	(in == 8'h69) ? 12'h2b6 : 
	(in == 8'h6a) ? 12'h2c4 : 
	(in == 8'h6b) ? 12'h2d1 : 
	(in == 8'h6c) ? 12'h2df : 
	(in == 8'h6d) ? 12'h2ec : 
	(in == 8'h6e) ? 12'h2fa : 
	(in == 8'h6f) ? 12'h308 : 
	(in == 8'h70) ? 12'h316 : 
	(in == 8'h71) ? 12'h324 : 
	(in == 8'h72) ? 12'h332 : 
	(in == 8'h73) ? 12'h341 : 
	(in == 8'h74) ? 12'h34f : 
	(in == 8'h75) ? 12'h35e : 
	(in == 8'h76) ? 12'h36d : 
	(in == 8'h77) ? 12'h37c : 
	(in == 8'h78) ? 12'h38b : 
	(in == 8'h79) ? 12'h39a : 
	(in == 8'h7a) ? 12'h3a9 : 
	(in == 8'h7b) ? 12'h3b9 : 
	(in == 8'h7c) ? 12'h3c8 : 
	(in == 8'h7d) ? 12'h3d8 : 
	(in == 8'h7e) ? 12'h3e8 : 
	(in == 8'h7f) ? 12'h3f8 : 
	(in == 8'h80) ? 12'h408 : 
	(in == 8'h81) ? 12'h418 : 
	(in == 8'h82) ? 12'h428 : 
	(in == 8'h83) ? 12'h439 : 
	(in == 8'h84) ? 12'h449 : 
	(in == 8'h85) ? 12'h45a : 
	(in == 8'h86) ? 12'h46b : 
	(in == 8'h87) ? 12'h47c : 
	(in == 8'h88) ? 12'h48d : 
	(in == 8'h89) ? 12'h49e : 
	(in == 8'h8a) ? 12'h4af : 
	(in == 8'h8b) ? 12'h4c1 : 
	(in == 8'h8c) ? 12'h4d2 : 
	(in == 8'h8d) ? 12'h4e4 : 
	(in == 8'h8e) ? 12'h4f6 : 
	(in == 8'h8f) ? 12'h508 : 
	(in == 8'h90) ? 12'h51a : 
	(in == 8'h91) ? 12'h52c : 
	(in == 8'h92) ? 12'h53e : 
	(in == 8'h93) ? 12'h551 : 
	(in == 8'h94) ? 12'h563 : 
	(in == 8'h95) ? 12'h576 : 
	(in == 8'h96) ? 12'h589 : 
	(in == 8'h97) ? 12'h59c : 
	(in == 8'h98) ? 12'h5af : 
	(in == 8'h99) ? 12'h5c2 : 
	(in == 8'h9a) ? 12'h5d6 : 
	(in == 8'h9b) ? 12'h5e9 : 
	(in == 8'h9c) ? 12'h5fd : 
	(in == 8'h9d) ? 12'h610 : 
	(in == 8'h9e) ? 12'h624 : 
	(in == 8'h9f) ? 12'h638 : 
	(in == 8'ha0) ? 12'h64c : 
	(in == 8'ha1) ? 12'h660 : 
	(in == 8'ha2) ? 12'h675 : 
	(in == 8'ha3) ? 12'h689 : 
	(in == 8'ha4) ? 12'h69e : 
	(in == 8'ha5) ? 12'h6b3 : 
	(in == 8'ha6) ? 12'h6c7 : 
	(in == 8'ha7) ? 12'h6dc : 
	(in == 8'ha8) ? 12'h6f1 : 
	(in == 8'ha9) ? 12'h707 : 
	(in == 8'haa) ? 12'h71c : 
	(in == 8'hab) ? 12'h731 : 
	(in == 8'hac) ? 12'h747 : 
	(in == 8'had) ? 12'h75d : 
	(in == 8'hae) ? 12'h773 : 
	(in == 8'haf) ? 12'h789 : 
	(in == 8'hb0) ? 12'h79f : 
	(in == 8'hb1) ? 12'h7b5 : 
	(in == 8'hb2) ? 12'h7cb : 
	(in == 8'hb3) ? 12'h7e2 : 
	(in == 8'hb4) ? 12'h7f8 : 
	(in == 8'hb5) ? 12'h80f : 
	(in == 8'hb6) ? 12'h826 : 
	(in == 8'hb7) ? 12'h83d : 
	(in == 8'hb8) ? 12'h854 : 
	(in == 8'hb9) ? 12'h86b : 
	(in == 8'hba) ? 12'h883 : 
	(in == 8'hbb) ? 12'h89a : 
	(in == 8'hbc) ? 12'h8b2 : 
	(in == 8'hbd) ? 12'h8ca : 
	(in == 8'hbe) ? 12'h8e1 : 
	(in == 8'hbf) ? 12'h8f9 : 
	(in == 8'hc0) ? 12'h912 : 
	(in == 8'hc1) ? 12'h92a : 
	(in == 8'hc2) ? 12'h942 : 
	(in == 8'hc3) ? 12'h95b : 
	(in == 8'hc4) ? 12'h973 : 
	(in == 8'hc5) ? 12'h98c : 
	(in == 8'hc6) ? 12'h9a5 : 
	(in == 8'hc7) ? 12'h9be : 
	(in == 8'hc8) ? 12'h9d7 : 
	(in == 8'hc9) ? 12'h9f0 : 
	(in == 8'hca) ? 12'ha0a : 
	(in == 8'hcb) ? 12'ha23 : 
	(in == 8'hcc) ? 12'ha3d : 
	(in == 8'hcd) ? 12'ha57 : 
	(in == 8'hce) ? 12'ha70 : 
	(in == 8'hcf) ? 12'ha8a : 
	(in == 8'hd0) ? 12'haa5 : 
	(in == 8'hd1) ? 12'habf : 
	(in == 8'hd2) ? 12'had9 : 
	(in == 8'hd3) ? 12'haf4 : 
	(in == 8'hd4) ? 12'hb0e : 
	(in == 8'hd5) ? 12'hb29 : 
	(in == 8'hd6) ? 12'hb44 : 
	(in == 8'hd7) ? 12'hb5f : 
	(in == 8'hd8) ? 12'hb7a : 
	(in == 8'hd9) ? 12'hb95 : 
	(in == 8'hda) ? 12'hbb1 : 
	(in == 8'hdb) ? 12'hbcc : 
	(in == 8'hdc) ? 12'hbe8 : 
	(in == 8'hdd) ? 12'hc04 : 
	(in == 8'hde) ? 12'hc20 : 
	(in == 8'hdf) ? 12'hc3c : 
	(in == 8'he0) ? 12'hc58 : 
	(in == 8'he1) ? 12'hc74 : 
	(in == 8'he2) ? 12'hc91 : 
	(in == 8'he3) ? 12'hcad : 
	(in == 8'he4) ? 12'hcca : 
	(in == 8'he5) ? 12'hce7 : 
	(in == 8'he6) ? 12'hd03 : 
	(in == 8'he7) ? 12'hd20 : 
	(in == 8'he8) ? 12'hd3e : 
	(in == 8'he9) ? 12'hd5b : 
	(in == 8'hea) ? 12'hd78 : 
	(in == 8'heb) ? 12'hd96 : 
	(in == 8'hec) ? 12'hdb3 : 
	(in == 8'hed) ? 12'hdd1 : 
	(in == 8'hee) ? 12'hdef : 
	(in == 8'hef) ? 12'he0d : 
	(in == 8'hf0) ? 12'he2b : 
	(in == 8'hf1) ? 12'he4a : 
	(in == 8'hf2) ? 12'he68 : 
	(in == 8'hf3) ? 12'he87 : 
	(in == 8'hf4) ? 12'hea5 : 
	(in == 8'hf5) ? 12'hec4 : 
	(in == 8'hf6) ? 12'hee3 : 
	(in == 8'hf7) ? 12'hf02 : 
	(in == 8'hf8) ? 12'hf21 : 
	(in == 8'hf9) ? 12'hf41 : 
	(in == 8'hfa) ? 12'hf60 : 
	(in == 8'hfb) ? 12'hf80 : 
	(in == 8'hfc) ? 12'hf9f : 
	(in == 8'hfd) ? 12'hfbf : 
	(in == 8'hfe) ? 12'hfdf : 
	12'h0ff;
endmodule
