module gamma(input [7:0] in, output reg [11:0] out);
always @(in) begin
case(in)
	8'h00: out = 12'h000;
	8'h01: out = 12'h000;
	8'h02: out = 12'h000;
	8'h03: out = 12'h000;
	8'h04: out = 12'h000;
	8'h05: out = 12'h000;
	8'h06: out = 12'h000;
	8'h07: out = 12'h000;
	8'h08: out = 12'h000;
	8'h09: out = 12'h000;
	8'h0a: out = 12'h000;
	8'h0b: out = 12'h000;
	8'h0c: out = 12'h000;
	8'h0d: out = 12'h000;
	8'h0e: out = 12'h000;
	8'h0f: out = 12'h000;
	8'h10: out = 12'h000;
	8'h11: out = 12'h000;
	8'h12: out = 12'h000;
	8'h13: out = 12'h000;
	8'h14: out = 12'h000;
	8'h15: out = 12'h000;
	8'h16: out = 12'h000;
	8'h17: out = 12'h000;
	8'h18: out = 12'h000;
	8'h19: out = 12'h000;
	8'h1a: out = 12'h000;
	8'h1b: out = 12'h001;
	8'h1c: out = 12'h001;
	8'h1d: out = 12'h001;
	8'h1e: out = 12'h001;
	8'h1f: out = 12'h001;
	8'h20: out = 12'h001;
	8'h21: out = 12'h001;
	8'h22: out = 12'h001;
	8'h23: out = 12'h001;
	8'h24: out = 12'h002;
	8'h25: out = 12'h002;
	8'h26: out = 12'h002;
	8'h27: out = 12'h002;
	8'h28: out = 12'h002;
	8'h29: out = 12'h003;
	8'h2a: out = 12'h003;
	8'h2b: out = 12'h003;
	8'h2c: out = 12'h004;
	8'h2d: out = 12'h004;
	8'h2e: out = 12'h004;
	8'h2f: out = 12'h005;
	8'h30: out = 12'h005;
	8'h31: out = 12'h006;
	8'h32: out = 12'h006;
	8'h33: out = 12'h007;
	8'h34: out = 12'h007;
	8'h35: out = 12'h008;
	8'h36: out = 12'h008;
	8'h37: out = 12'h009;
	8'h38: out = 12'h00a;
	8'h39: out = 12'h00a;
	8'h3a: out = 12'h00b;
	8'h3b: out = 12'h00c;
	8'h3c: out = 12'h00d;
	8'h3d: out = 12'h00d;
	8'h3e: out = 12'h00e;
	8'h3f: out = 12'h00f;
	8'h40: out = 12'h010;
	8'h41: out = 12'h011;
	8'h42: out = 12'h012;
	8'h43: out = 12'h014;
	8'h44: out = 12'h015;
	8'h45: out = 12'h016;
	8'h46: out = 12'h017;
	8'h47: out = 12'h019;
	8'h48: out = 12'h01a;
	8'h49: out = 12'h01c;
	8'h4a: out = 12'h01d;
	8'h4b: out = 12'h01f;
	8'h4c: out = 12'h020;
	8'h4d: out = 12'h022;
	8'h4e: out = 12'h024;
	8'h4f: out = 12'h026;
	8'h50: out = 12'h028;
	8'h51: out = 12'h02a;
	8'h52: out = 12'h02c;
	8'h53: out = 12'h02e;
	8'h54: out = 12'h030;
	8'h55: out = 12'h033;
	8'h56: out = 12'h035;
	8'h57: out = 12'h037;
	8'h58: out = 12'h03a;
	8'h59: out = 12'h03d;
	8'h5a: out = 12'h040;
	8'h5b: out = 12'h042;
	8'h5c: out = 12'h045;
	8'h5d: out = 12'h048;
	8'h5e: out = 12'h04c;
	8'h5f: out = 12'h04f;
	8'h60: out = 12'h052;
	8'h61: out = 12'h056;
	8'h62: out = 12'h059;
	8'h63: out = 12'h05d;
	8'h64: out = 12'h061;
	8'h65: out = 12'h065;
	8'h66: out = 12'h069;
	8'h67: out = 12'h06d;
	8'h68: out = 12'h071;
	8'h69: out = 12'h076;
	8'h6a: out = 12'h07a;
	8'h6b: out = 12'h07f;
	8'h6c: out = 12'h084;
	8'h6d: out = 12'h089;
	8'h6e: out = 12'h08e;
	8'h6f: out = 12'h093;
	8'h70: out = 12'h098;
	8'h71: out = 12'h09e;
	8'h72: out = 12'h0a4;
	8'h73: out = 12'h0a9;
	8'h74: out = 12'h0af;
	8'h75: out = 12'h0b5;
	8'h76: out = 12'h0bc;
	8'h77: out = 12'h0c2;
	8'h78: out = 12'h0c9;
	8'h79: out = 12'h0d0;
	8'h7a: out = 12'h0d7;
	8'h7b: out = 12'h0de;
	8'h7c: out = 12'h0e5;
	8'h7d: out = 12'h0ec;
	8'h7e: out = 12'h0f4;
	8'h7f: out = 12'h0fc;
	8'h80: out = 12'h104;
	8'h81: out = 12'h10c;
	8'h82: out = 12'h115;
	8'h83: out = 12'h11d;
	8'h84: out = 12'h126;
	8'h85: out = 12'h12f;
	8'h86: out = 12'h138;
	8'h87: out = 12'h142;
	8'h88: out = 12'h14b;
	8'h89: out = 12'h155;
	8'h8a: out = 12'h15f;
	8'h8b: out = 12'h16a;
	8'h8c: out = 12'h174;
	8'h8d: out = 12'h17f;
	8'h8e: out = 12'h18a;
	8'h8f: out = 12'h195;
	8'h90: out = 12'h1a0;
	8'h91: out = 12'h1ac;
	8'h92: out = 12'h1b8;
	8'h93: out = 12'h1c4;
	8'h94: out = 12'h1d1;
	8'h95: out = 12'h1dd;
	8'h96: out = 12'h1ea;
	8'h97: out = 12'h1f8;
	8'h98: out = 12'h205;
	8'h99: out = 12'h213;
	8'h9a: out = 12'h221;
	8'h9b: out = 12'h22f;
	8'h9c: out = 12'h23e;
	8'h9d: out = 12'h24c;
	8'h9e: out = 12'h25c;
	8'h9f: out = 12'h26b;
	8'ha0: out = 12'h27b;
	8'ha1: out = 12'h28b;
	8'ha2: out = 12'h29b;
	8'ha3: out = 12'h2ac;
	8'ha4: out = 12'h2bd;
	8'ha5: out = 12'h2ce;
	8'ha6: out = 12'h2df;
	8'ha7: out = 12'h2f1;
	8'ha8: out = 12'h303;
	8'ha9: out = 12'h316;
	8'haa: out = 12'h329;
	8'hab: out = 12'h33c;
	8'hac: out = 12'h350;
	8'had: out = 12'h364;
	8'hae: out = 12'h378;
	8'haf: out = 12'h38c;
	8'hb0: out = 12'h3a1;
	8'hb1: out = 12'h3b7;
	8'hb2: out = 12'h3cc;
	8'hb3: out = 12'h3e2;
	8'hb4: out = 12'h3f9;
	8'hb5: out = 12'h40f;
	8'hb6: out = 12'h427;
	8'hb7: out = 12'h43e;
	8'hb8: out = 12'h456;
	8'hb9: out = 12'h46e;
	8'hba: out = 12'h487;
	8'hbb: out = 12'h4a0;
	8'hbc: out = 12'h4ba;
	8'hbd: out = 12'h4d4;
	8'hbe: out = 12'h4ee;
	8'hbf: out = 12'h509;
	8'hc0: out = 12'h524;
	8'hc1: out = 12'h540;
	8'hc2: out = 12'h55c;
	8'hc3: out = 12'h578;
	8'hc4: out = 12'h595;
	8'hc5: out = 12'h5b3;
	8'hc6: out = 12'h5d1;
	8'hc7: out = 12'h5ef;
	8'hc8: out = 12'h60e;
	8'hc9: out = 12'h62d;
	8'hca: out = 12'h64c;
	8'hcb: out = 12'h66d;
	8'hcc: out = 12'h68d;
	8'hcd: out = 12'h6ae;
	8'hce: out = 12'h6d0;
	8'hcf: out = 12'h6f2;
	8'hd0: out = 12'h715;
	8'hd1: out = 12'h738;
	8'hd2: out = 12'h75c;
	8'hd3: out = 12'h780;
	8'hd4: out = 12'h7a4;
	8'hd5: out = 12'h7c9;
	8'hd6: out = 12'h7ef;
	8'hd7: out = 12'h815;
	8'hd8: out = 12'h83c;
	8'hd9: out = 12'h863;
	8'hda: out = 12'h88b;
	8'hdb: out = 12'h8b4;
	8'hdc: out = 12'h8dd;
	8'hdd: out = 12'h906;
	8'hde: out = 12'h930;
	8'hdf: out = 12'h95b;
	8'he0: out = 12'h986;
	8'he1: out = 12'h9b2;
	8'he2: out = 12'h9df;
	8'he3: out = 12'ha0c;
	8'he4: out = 12'ha39;
	8'he5: out = 12'ha67;
	8'he6: out = 12'ha96;
	8'he7: out = 12'hac6;
	8'he8: out = 12'haf6;
	8'he9: out = 12'hb26;
	8'hea: out = 12'hb58;
	8'heb: out = 12'hb8a;
	8'hec: out = 12'hbbc;
	8'hed: out = 12'hbf0;
	8'hee: out = 12'hc23;
	8'hef: out = 12'hc58;
	8'hf0: out = 12'hc8d;
	8'hf1: out = 12'hcc3;
	8'hf2: out = 12'hcfa;
	8'hf3: out = 12'hd31;
	8'hf4: out = 12'hd69;
	8'hf5: out = 12'hda1;
	8'hf6: out = 12'hddb;
	8'hf7: out = 12'he15;
	8'hf8: out = 12'he50;
	8'hf9: out = 12'he8b;
	8'hfa: out = 12'hec7;
	8'hfb: out = 12'hf04;
	8'hfc: out = 12'hf42;
	8'hfd: out = 12'hf80;
	8'hfe: out = 12'hfbf;
	8'hff: out = 12'hfff;
endcase
end
endmodule
